module LOBA_LOB_16 (x, y);
    input [15:0] x;
    output reg [15:0] y;

    always @ (*) begin
        if (x[15])
            y <= 16'b1000000000000000;
        else if (x[14])
            y <= 16'b0100000000000000;
        else if (x[13])
            y <= 16'b0010000000000000;
        else if (x[12])
            y <= 16'b0001000000000000;
        else if (x[11])
            y <= 16'b0000100000000000;
        else if (x[10])
            y <= 16'b0000010000000000;
        else if (x[9])
            y <= 16'b0000001000000000;
        else if (x[8])
            y <= 16'b0000000100000000;
        else if (x[7])
            y <= 16'b0000000010000000;
        else if (x[6])
            y <= 16'b0000000001000000;
        else if (x[5])
            y <= 16'b0000000000100000;
        else if (x[4])
            y <= 16'b0000000000010000;
        else if (x[3])
            y <= 16'b0000000000001000;
        else if (x[2])
            y <= 16'b0000000000000100;
        else if (x[1])
            y <= 16'b0000000000000010;
        else if (x[0])
            y <= 16'b0000000000000001;
        else
            y <= 16'b0000000000000000;
    end
endmodule
